<?xml version="1.0" encoding="utf-8"?>
<!-- Generator: Adobe Illustrator 17.0.0, SVG Export Plug-In . SVG Version: 6.00 Build 0)  -->
<!DOCTYPE svg PUBLIC "-//W3C//DTD SVG 1.1//EN" "http://www.w3.org/Graphics/SVG/1.1/DTD/svg11.dtd">
<svg version="1.1" id="Layer_1" xmlns="http://www.w3.org/2000/svg" xmlns:xlink="http://www.w3.org/1999/xlink" x="0px" y="0px"
	 width="203px" height="72.737px" viewBox="422.667 409.934 203 72.737" enable-background="new 422.667 409.934 203 72.737"
	 xml:space="preserve">
<linearGradient id="SVGID_1_" gradientUnits="userSpaceOnUse" x1="443.667" y1="557.12" x2="610.3448" y2="557.12" gradientTransform="matrix(1 0 0 -1 -21 1003.5)">
	<stop  offset="0" style="stop-color:#F7941E"/>
	<stop  offset="0.2135" style="stop-color:#F3961F"/>
	<stop  offset="0.404" style="stop-color:#E99B22"/>
	<stop  offset="0.5857" style="stop-color:#D6A328"/>
	<stop  offset="0.762" style="stop-color:#BDAF30"/>
	<stop  offset="0.9329" style="stop-color:#9CBF3A"/>
	<stop  offset="1" style="stop-color:#8DC63F"/>
</linearGradient>
<path fill="url(#SVGID_1_)" d="M592.235,440.833c-1.721-5.047-5.086-7.571-10.096-7.571c0,0-4.291,0-4.361,0
	c-0.07,0-0.113,0.059-0.113,0.204c0,1.103,0.478,2.032,1.432,2.697c0.159,0.111,0.4,0.353,1.12,0.353
	c2.567,0,4.223,0.051,6.222,1.546c1.868,1.397,2.813,3.687,2.813,6.902v34.191c0,2.448,1.103,3.671,3.328,3.671
	c0.138,0,0.229-0.124,0.229-0.23s0-37.287,0-37.287C592.809,443.74,592.619,442.248,592.235,440.833z M535.988,467.34
	c0.135,0,17.022,0,17.022,0c2.255,0,3.382-1.315,3.382-3.945v-1.803c0-2.311-0.3-4.227-0.902-5.749
	c-1.634-4.358-5.053-6.538-10.891-6.538c-5.148,0-7.191,1.386-8.612,2.572c-2.404,2.005-3.606,5.055-3.606,9.152v11.611l0.226,2.03
	c1.259,5.336,5.053,8.003,11.385,8.003c0,0,12.106,0,12.175,0c0.172,0,0.225-0.112,0.185-0.273c-0.015-0.06-0.11-0.678-0.298-1.193
	c-0.469-1.283-1.691-1.916-3.72-1.916c0,0-4.124,0-6.426,0c-2.301,0-4.217-0.012-5.186-0.338c-3.304-1.114-4.959-3.4-4.959-6.876
	c0,0,0-4.424,0-4.509C535.763,467.48,535.853,467.34,535.988,467.34z M535.763,462.268c0-2.292,0.149-4.02,0.45-5.185
	c1.051-2.932,3.721-4.397,8.398-4.397c5.904,0,8.399,2.818,8.399,8.454v1.24c0,1.128-0.564,1.691-1.691,1.691h-15.556V462.268z
	 M519.088,438.108c-1.29,1.82-1.934,4.124-1.934,6.912c0,0,0,33.519,0,33.916c0,0.767,0.202,1.374,0.385,1.823
	c0.52,1.275,1.483,1.912,2.885,1.912c0.109,0,0.225-0.045,0.225-0.225c0-0.179,0-26.604,0-26.604s3.786,0,5.752,0
	c2.225,0,3.605-1.14,3.605-2.931c0-0.225-0.075-0.338-0.225-0.338h-9.131c0,0,0-6.919,0-7.44s0.188-2.211,0.297-2.604
	c0.922-3.338,3.066-5.173,6.017-5.173c3.381-0.263,5.072-1.278,5.072-3.044c0-0.372,0-0.451-0.259-0.451c-0.828,0-3.383,0-3.919,0
	C522.943,433.86,520.327,436.358,519.088,438.108z M495.778,449.191c-0.119,0-12.799,0-13.464,0c-0.887,0-2.205,0.226-2.205,0.226
	c-5.487,1.26-8.229,4.791-8.229,10.596c0,0,0,22.324,0,22.434s0.093,0.225,0.226,0.225c0.092,0,11.836,0,11.836,0
	c3.926,0,6.782-0.939,8.568-2.818h0.112c0,1.56,1.014,2.499,3.044,2.818c0.225,0,0.338-0.074,0.338-0.225c0,0,0-32.911,0-33.03
	C496.004,449.299,495.897,449.191,495.778,449.191z M492.509,470.835c0,1.109-0.19,2.751-0.451,3.607
	c-0.261,0.856-1.153,2.176-2,2.92c-1.376,1.21-3.227,1.814-5.553,1.814h-9.019c0,0,0-18.731,0-19.502
	c0-0.771,0.127-1.766,0.339-2.592c0.245-0.954,1.285-2.323,2.248-3.041c1.223-0.913,2.796-1.356,4.74-1.356h9.695V470.835
	L492.509,470.835z M510.441,449.417c-2.828,0-4.566,0.826-6.539,2.479h-0.112c0-1.115-0.851-1.926-2.553-2.434
	c-0.19-0.057-0.457-0.135-0.603-0.159c-0.114-0.019-0.226,0.07-0.226,0.225s0,29.294,0,29.648c0,0.463-0.043,0.856,0.113,1.241
	c0.63,1.549,1.619,2.254,3.156,2.254c0.187,0,0.225-0.138,0.225-0.225s0-21.643,0-21.643c0-2.099,0.577-3.928,1.254-5.104
	c0.796-1.382,3.141-3.013,4.674-3.013c1.559,0,2.504-0.9,2.928-2.701c0.018-0.075,0.05-0.258,0.05-0.344s-0.073-0.225-0.225-0.225
	C512.43,449.417,510.441,449.417,510.441,449.417z M455.923,449.303h-1.24c-4.454,0-7.609,1.504-9.47,4.509h-0.337
	c-1.861-3.006-4.943-4.509-9.244-4.509h-2.48c-2.762,0-5.129,0.902-7.102,2.705c-0.282-1.803-1.319-2.705-3.156-2.705
	c-0.126,0-0.226,0.142-0.226,0.225c0,0.083,0,29.838,0,30.009c0,0.531,0.166,0.805,0.262,1.024c0.615,1.406,1.584,2.109,2.896,2.109
	c0.113,0,0.225-0.102,0.225-0.225c0-0.123,0-21.982,0-21.982c0-1.033,0.188-2.199,0.563-3.495c1.298-2.856,3.626-4.284,6.991-4.284
	h2.141c1.145,0,2.385,0.262,3.719,0.789c2.555,1.184,3.833,3.739,3.833,7.665c0,0,0,18.179,0,18.375
	c0,0.197,0.113,0.675,0.113,0.675c0.526,1.654,1.524,2.48,3.044,2.48c0.109,0,0.225-0.08,0.225-0.225c0-0.145,0-20.518,0-20.518
	c0-2.629,0.3-4.508,0.902-5.635c1.127-2.405,3.458-3.607,6.99-3.607h1.578c5.26,0,7.892,3.156,7.892,9.469c0,0,0,16.766,0,16.905
	c0,0.366,0.041,0.529,0.067,0.671c0.354,1.961,1.346,2.94,2.976,2.94c0.225,0,0.338-0.074,0.338-0.225v-20.855
	c0-2.988-0.489-5.28-1.466-6.877C464.264,451.108,460.919,449.303,455.923,449.303z M625.358,409.935c-0.127,0-15.05,0-15.05,0
	v-0.001c0,0-0.949,0-6.712,0s-9.336,2.743-10.596,8.229c0,0-0.225,1.385-0.225,1.917s0,13.468,0,13.538
	c0,0.335,0.091,0.44,0.415,0.44c0.134,0,14.945,0,14.945,0v0.001h6.712c5.805,0,9.336-2.743,10.596-8.229
	c0,0,0.225-0.999,0.225-1.917s0-13.578,0-13.69C625.667,410.11,625.561,409.935,625.358,409.935z M622.172,423.125
	c0,3.476-1.398,5.77-4.397,6.988c-0.495,0.201-1.889,0.451-4.255,0.451s-17.252,0-17.252,0v-9.695c0-3.476,1.418-5.751,4.397-6.988
	c0.835-0.347,1.772-0.339,2.592-0.339s5.342,0,5.342,0c0,0.001,0,0.001,0,0.002h13.574V423.125z M564.271,467.34
	c0.135,0,17.022,0,17.022,0c2.255,0,3.382-1.315,3.382-3.945v-1.803c0-2.311-0.3-4.227-0.902-5.749
	c-1.634-4.358-5.053-6.538-10.891-6.538c-5.148,0-7.191,1.386-8.612,2.572c-2.404,2.005-3.606,5.055-3.606,9.152v11.611l0.226,2.03
	c1.259,5.336,5.053,8.003,11.385,8.003c0,0,12.106,0,12.175,0c0.172,0,0.225-0.112,0.185-0.273c-0.015-0.06-0.11-0.678-0.298-1.193
	c-0.469-1.283-1.691-1.916-3.72-1.916c0,0-4.125,0-6.426,0c-2.301,0-4.217-0.012-5.186-0.338c-3.304-1.114-4.959-3.4-4.959-6.876
	c0,0,0-4.424,0-4.509C564.046,467.48,564.135,467.34,564.271,467.34z M564.046,462.268c0-2.292,0.149-4.02,0.45-5.185
	c1.051-2.932,3.721-4.397,8.398-4.397c5.904,0,8.399,2.818,8.399,8.454v1.24c0,1.128-0.564,1.691-1.691,1.691h-15.556V462.268z"/>
</svg>
